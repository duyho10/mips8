module Nor_1bit(c,a,b);
input a,b;
output c;
nor (c,a,b);
endmodule
