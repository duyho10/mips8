module Or_1bit(c,a,b);
input a,b;
output c;
or (c,a,b);
endmodule
