module And_1bit(c,a,b);
input a,b;
output c;
and (c,a,b);
endmodule
