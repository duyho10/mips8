module Xor_1bit(c,a,b);
input a,b;
output c;
xor (c,a,b);
endmodule
